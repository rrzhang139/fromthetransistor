module mux4 (
    input wire [1:0] sel,  // 2-bit select signal
    input wire [3:0] in,   // 4-bit input data
    output wire out        // Output data
);

    always @(sel, in) begin
        case(sel)
            2'b00: out = in[0];
            2'b01: out = in[1];
            2'b10: out = in[2];
            2'b11: out = in[3];
        endcase
    end

endmodule
